LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_TEXTIO.all;
use STD.TEXTIO.all;

USE WORK.UTILITIES.ALL;

ENTITY TESTBENCH IS
END ENTITY;

ARCHITECTURE BEHAVIOUR OF TESTBENCH IS

COMPONENT IITBProc is
	port( 
		clk, load: in std_logic;
		DataIn: in std_logic_vector (15 downto 0);
		Interface: out d2;
		Trap: out std_logic);
END COMPONENT;

SIGNAL CLK, LOAD, TRAP: STD_LOGIC;
SIGNAL DATAIN: STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL INTERFACE: d2;

BEGIN

	CPU_INST: IITBProc
		PORT MAP (CLK, LOAD, DATAIN, INTERFACE, TRAP);
	
	PROCESS
		FILE INPUT_FILE: TEXT OPEN READ_MODE IS "/home/burixzura/acads/CS 254/Project/GitHub/IITB-Proc/instructions/jlr1.txt";
		VARIABLE INPUT_LINE: LINE;
		VARIABLE INPUT_VAR: STD_LOGIC_VECTOR (15 DOWNTO 0);
		VARIABLE INIT: STD_LOGIC := '0';
	BEGIN
	
		
		IF (INIT='0') THEN
			LOAD <= '1';
			FOR I IN 0 TO 1 LOOP
				IF (I=0) THEN
					WHILE NOT ENDFILE(INPUT_FILE) LOOP
						CLK <= '0';
						WAIT FOR 50 NS;
						CLK <= '1';
						READLINE(INPUT_FILE, INPUT_LINE);
						READ(INPUT_LINE, INPUT_VAR);
						DATAIN <= INPUT_VAR;
						WAIT FOR 50 NS;
					END LOOP;
				ELSE
					CLK <= '0';
					WAIT FOR 50 NS;
					CLK <= '1';
					DATAIN <= "1111111111111111";
					WAIT FOR 50 NS;
				END IF;
			END LOOP;
			INIT:='1';
		ELSE
			LOAD <= '0';
			CLK <= '0';
			WAIT FOR 50 NS;
			CLK <= '1';
			WAIT FOR 50 NS;
			IF (TRAP='1') THEN
				WAIT;
			END IF;
		END IF;
		
	END PROCESS;

END ARCHITECTURE;
