library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package utilities is

	type d2 is array (0 to 7) of std_logic_vector (15 downto 0);

end package;