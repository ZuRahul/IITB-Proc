LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TESTBENCH IS
END ENTITY;

ARCHITECTURE BEHAVIOUR OF TESTBENCH IS

COMPONENT IITBProc is
	port( 
		clk, load: in std_logic;
		DataIn: in std_logic_vector (15 downto 0));
END COMPONENT;

SIGNAL CLK, LOAD: STD_LOGIC;
SIGNAL DATAIN: STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN

	CPU_INST: IITBProc
		PORT MAP (CLK, LOAD, DATAIN);
	
	PROCESS
		FILE INPUT_FILE: TEXT OPEN READ_MODE IS "instructions.txt";
		VARIABLE INPUT_LINE: LINE;
		VARIABLE INPUT_VAR: STD_LOGIC_VECTOR (15 DOWNTO 0);
	BEGIN
	
		FOR I IN 0 TO 1 LOOP
		 IF (I=0) THEN
			LOAD <= '1';
			WHILE NOT ENDFILE(INPUT_FILE) LOOP
				CLK <= '0';
				WAIT FOR 10 NS;
				CLK<='1';
				READLINE(INPUT_FILE, INPUT_LINE);
				READ(INPUT_LINE, INPUT_VAR);
				DATAIN <= INPUT_VAR;
				WAIT FOR 10 NS;
			END LOOP;
		 ELSE
			LOAD <= '0';
			
		 END IF;
		END LOOP;
	END PROCESS;

END ARCHITECTURE;